module f_adder(A,B,op);
input [15:0] A,B;
output [15:0] op;
reg sign;
reg [4:0] exp;
reg [9:0] man;


endmodule