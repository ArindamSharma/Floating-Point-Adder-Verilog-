module f_adder(A,B)

endmodule