module f_adder(A,B,op);
input [15:0] A,B;
output [15:0] op;
reg sign;
reg [0:4] exp;
reg [0:9] man;


endmodule